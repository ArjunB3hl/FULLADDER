* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT efuse PLUS MINUS
.ENDS
***************************************
.SUBCKT hvpwdnwhvnw_dio_hvpw_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT lcesd1_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT lcesd2_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT lowcpad_rf APAD AVSS
.ENDS
***************************************
.SUBCKT lvpwdnwhvnw_dio_hvpw_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin_hl TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_1p0_sin_hl_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_1p5_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_1p5_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_shield PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3ds TOP BOTTOM
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3ds_3t TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_wos PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_4p0_sin_3dshs TOP BOTTOM
.ENDS
***************************************
.SUBCKT mimcap_4p0_sin_3dshs_3t TOP BOTTOM GNODE
.ENDS
***************************************
.SUBCKT mimcap_shield PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_wos PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nch_hv5_5vnw_ac D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT nch_hva_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hva_ndd_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvau_ndd_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvi_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nch_hviah_ndd_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvish_nbl_mac D G S B NBL_ISO SUB
.ENDS
***************************************
.SUBCKT nch_hvish_ndd_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvisl_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvnw_6t D G S B HVNW_ISO SUB
.ENDS
***************************************
.SUBCKT nch_hvs_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvs_ndd_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvsl_mac D G S B
.ENDS
***************************************
.SUBCKT nch_hvsu_ndd_mac D G S B
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT ndio_sbd_mac PLUS MINUS
.ENDS
***************************************
.SUBCKT ndld24_g5_ac D G BS SUB
.ENDS
***************************************
.SUBCKT ndld40_g5_ac D G BS SUB
.ENDS
***************************************
.SUBCKT nhvpwdnw10_4t C B E SUB
.ENDS
***************************************
.SUBCKT nhvpwdnw5_4t C B E SUB
.ENDS
***************************************
.SUBCKT nld12_g12_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld12_g2_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld14_g12_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld14_g2_mac D G BS SUB
.ENDS
***************************************
.SUBCKT nld18_g5_ac D G BS SUB
.ENDS
***************************************
.SUBCKT nld24_g5_ac D G BS SUB
.ENDS
***************************************
.SUBCKT nld32_g5_ac D G BS SUB
.ENDS
***************************************
.SUBCKT nld40_g5_ac D G BS SUB
.ENDS
***************************************
.SUBCKT nld60_g5_ac D G BS SUB
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33_mis PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_mis PLUS MINUS
.ENDS
***************************************
.SUBCKT nvmrpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT pa18_g5_ac D G S B SUB
.ENDS
***************************************
.SUBCKT pa24_g5_ac D G S B SUB
.ENDS
***************************************
.SUBCKT pa32_g5_ac D G S B SUB
.ENDS
***************************************
.SUBCKT pa40_g5_full_soa_ac D G S B SUB
.ENDS
***************************************
.SUBCKT pa40_g5_low_ron_ac D G S B SUB
.ENDS
***************************************
.SUBCKT pa50_g5_ac D G S B SUB
.ENDS
***************************************
.SUBCKT pa60_g5_full_soa_ac D G S B SUB
.ENDS
***************************************
.SUBCKT pch_5t D G S B SUB
.ENDS
***************************************
.SUBCKT pch_hva_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pch_hva_pdd_mac D G S B
.ENDS
***************************************
.SUBCKT pch_hvau_pdd_mac D G S B
.ENDS
***************************************
.SUBCKT pch_hvs_mac D G S B SUB
.ENDS
***************************************
.SUBCKT pch_hvs_pdd_mac D G S B
.ENDS
***************************************
.SUBCKT pch_hvsl_mac D G S B
.ENDS
***************************************
.SUBCKT pch_hvsu_pdd_mac D G S B
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT phvnw_dio_hvpw_3t PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT rhim PLUS MINUS
.ENDS
***************************************
.SUBCKT rhvnw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rhvnw_60 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rhvnwhvpw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rhvpw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rhvpw_60 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rldpwod PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rldpwsti PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnddhvpw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_ell PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_ell_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_ull PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_ull_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_ell PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_ell_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_ull PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_ull_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpbody PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpddhvnw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpod_ell PLUS MINUS
.ENDS
***************************************
.SUBCKT rpod_ell_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_ull PLUS MINUS
.ENDS
***************************************
.SUBCKT rpod_ull_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_ell PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodrpo_ell_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_ull PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodrpo_ull_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_ell PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodw_ell_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_ull PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodw_ull_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri3k PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyhri3k_dis PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyhri_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_dio_60 PLUS MINUS
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nr36 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_w40 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT zd_dio_4t PLUS MINUS NBL_ISO SUB
.ENDS
***************************************
.SUBCKT PMOS 1 2 3 4
** N=5 EP=4 IP=0 FDC=2
M0 4 1 3 3 P L=1.8e-07 W=1e-06 $X=370 $Y=540 $D=39
M1 3 2 4 3 P L=1.8e-07 W=1e-06 $X=1100 $Y=540 $D=39
.ENDS
***************************************
.SUBCKT NMOS
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT FA A B C VSS VDD Co S
** N=23 EP=7 IP=25 FDC=36
M0 21 A VSS VSS N L=1.8e-07 W=1e-06 $X=3750 $Y=4910 $D=3
M1 3 B 21 VSS N L=1.8e-07 W=1e-06 $X=4480 $Y=4910 $D=3
M2 22 A VSS VSS N L=1.8e-07 W=1e-06 $X=6570 $Y=4910 $D=3
M3 4 3 22 VSS N L=1.8e-07 W=1e-06 $X=7300 $Y=4910 $D=3
M4 23 3 VSS VSS N L=1.8e-07 W=1e-06 $X=9390 $Y=4920 $D=3
M5 5 B 23 VSS N L=1.8e-07 W=1e-06 $X=10120 $Y=4920 $D=3
M6 15 4 VSS VSS N L=1.8e-07 W=2e-06 $X=12210 $Y=4910 $D=3
M7 7 5 15 VSS N L=1.8e-07 W=2e-06 $X=12940 $Y=4910 $D=3
M8 16 C VSS VSS N L=1.8e-07 W=4e-06 $X=15030 $Y=4910 $D=3
M9 8 7 16 VSS N L=1.8e-07 W=4e-06 $X=15760 $Y=4910 $D=3
M10 17 7 VSS VSS N L=1.8e-07 W=5e-06 $X=17850 $Y=4910 $D=3
M11 10 8 17 VSS N L=1.8e-07 W=5e-06 $X=18580 $Y=4910 $D=3
M12 18 8 VSS VSS N L=1.8e-07 W=5e-06 $X=20670 $Y=4910 $D=3
M13 9 C 18 VSS N L=1.8e-07 W=5e-06 $X=21400 $Y=4910 $D=3
M14 19 3 VSS VSS N L=1.8e-07 W=5e-06 $X=23490 $Y=4910 $D=3
M15 Co 8 19 VSS N L=1.8e-07 W=5e-06 $X=24220 $Y=4910 $D=3
M16 20 9 VSS VSS N L=1.8e-07 W=1.9e-05 $X=26310 $Y=4910 $D=3
M17 S 10 20 VSS N L=1.8e-07 W=1.9e-05 $X=27040 $Y=4910 $D=3
M18 5 3 VDD VDD P L=1.8e-07 W=1e-06 $X=9390 $Y=60720 $D=39
M19 VDD B 5 VDD P L=1.8e-07 W=1e-06 $X=10120 $Y=60720 $D=39
M20 7 4 VDD VDD P L=1.8e-07 W=2e-06 $X=12210 $Y=59710 $D=39
M21 VDD 5 7 VDD P L=1.8e-07 W=2e-06 $X=12940 $Y=59710 $D=39
M22 8 C VDD VDD P L=1.8e-07 W=4e-06 $X=15030 $Y=57710 $D=39
M23 VDD 7 8 VDD P L=1.8e-07 W=4e-06 $X=15760 $Y=57710 $D=39
M24 10 7 VDD VDD P L=1.8e-07 W=5e-06 $X=17850 $Y=56710 $D=39
M25 VDD 8 10 VDD P L=1.8e-07 W=5e-06 $X=18580 $Y=56710 $D=39
M26 9 8 VDD VDD P L=1.8e-07 W=5e-06 $X=20670 $Y=56710 $D=39
M27 VDD C 9 VDD P L=1.8e-07 W=5e-06 $X=21400 $Y=56710 $D=39
M28 Co 3 VDD VDD P L=1.8e-07 W=5e-06 $X=23490 $Y=56710 $D=39
M29 VDD 8 Co VDD P L=1.8e-07 W=5e-06 $X=24220 $Y=56710 $D=39
M30 S 9 VDD VDD P L=1.8e-07 W=1.9e-05 $X=26310 $Y=42710 $D=39
M31 VDD 10 S VDD P L=1.8e-07 W=1.9e-05 $X=27040 $Y=42710 $D=39
X32 A B VDD 3 PMOS $T=3380 60170 0 0 $X=2760 $Y=56910
X33 A 3 VDD 4 PMOS $T=6200 60170 0 0 $X=5580 $Y=56910
.ENDS
***************************************
